module nand_gate(input wire a, b, output wire out);
  assign out = ~(a & b);
endmodule